/home/arpit23132/Desktop/RISCV_Final/gsclib090_translated_ref.lef